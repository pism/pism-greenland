netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:output.checkpoint.interval = 48.0;
    
    pism_overrides:stress_balance.sia.max_diffusivity = 1000000.0;

    pism_overrides:surface.pdd.air_temp_all_precip_as_snow = 272.15;

    pism_overrides:surface.pdd.air_temp_all_precip_as_rain = 274.15;

    pism_overrides:surface.pdd.refreeze = 0.47;

    pism_overrides:surface.pdd.refreeze_ice_melt = "no";

    pism_overrides:run_info.institution = "University of Alaska Fairbanks";

    pism_overrides:surface.force_to_thickness.alpha = .8;

    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor = 1.0;

    pism_overrides:ocean.sub_shelf_heat_flux_into_ice = 50.0;

    pism_overrides:geometry.ice_free_thickness_standard = 10.0;

}
